LIBRARY IEEE;
USE IEEE.STD_logic_1164.ALL;
-----------------------------------------------------
ENTITY tb_Cnt4_e IS 
END tb_Cnt4_e;
-----------------------------------------
