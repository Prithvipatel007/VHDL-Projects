library IEEE;
USE IEEE.STD_LOGIC_1164.ALL;

ENTITY tb_txd_e IS 
END tb_txd_e;