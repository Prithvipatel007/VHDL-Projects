-- --------------------------------------------------------------------
-- --------------------------------------------------------------------
-- file: reg08_a1.vhd, last modified: 2021-1202
-- --------------------------------------------------------------------
-- --------------------------------------------------------------------
-- some GHDL-cmds:   ghdl -s xxx.vhd  : Syntax check
--                   ghdl -a xxx.vhd  : Assembles file xxx.vhd
--                   ghdl -e xyz      : Elaborates xyz
-- prepare waveform: ghdl -r xxx_TB1 --wave=xxx_TB1_wave.ghw
-- --------------------------------------------------------------------
-- --------------------------------------------------------------------
  LIBRARY IEEE;
  USE IEEE.STD_LOGIC_1164.ALL;
-- ------------------------------------------------------------
  ARCHITECTURE a1 OF reg08 IS

  SIGNAL st_s : STD_LOGIC_VECTOR (7 DOWNTO 0);
-- ------------------------------------------------------------
  BEGIN
  ldx : PROCESS (rb_i,cp_i,en_i,st_s)
   BEGIN
   IF (rb_i='0') THEN st_s <= X"00";
   ELSIF (cp_i='1' AND cp_i'EVENT)
    THEN
     IF  (en_i='1') THEN st_s(7 DOWNTO 0) <= d_i(7 DOWNTO 0);
     END IF;
   END IF;
   END PROCESS ldx;
-- ------------------------------------------------------------
  q_o(7 DOWNTO 0) <= st_s(7 DOWNTO 0);
-- ------------------------------------------------------------
  END a1;
-- ------------------------------------------------------------

