LIBRARY IEEE;
USE IEEE.std_logic_1164.ALL;
USE IEEE.numeric_std.ALL;

ENTITY sft_reg_tb IS
END sft_reg_tb;
-------------------------------------------------------------------