library ieee;
use ieee.std_logic_1164.all;

entity tb_baud_e is 
end tb_baud_e;

