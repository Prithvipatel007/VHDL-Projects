LIBRARY IEEE;
USE IEEE.STD_LOGIC_1164.ALL;
-----------------------------------------------------------
ENTITY tb_uart_ctrl_fsm_e IS 
END tb_uart_ctrl_fsm_e;

