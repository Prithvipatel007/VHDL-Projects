LIBRARY IEEE;
USE IEEE.STD_LOGIC_1164.ALL;

ENTITY tb_uart_tx_e IS
END tb_uart_tx_e;