-- --------------------------------------------------------------------
-- --------------------------------------------------------------------
-- file: uat_e.vhd, last modified: 2021-1208
-- --------------------------------------------------------------------
-- --------------------------------------------------------------------
  LIBRARY IEEE;
  USE IEEE.STD_LOGIC_1164.ALL;
--USE WORK.uat_pack.ALL;
-- --------------------------------------------------------------------
  ENTITY uat IS
   PORT (rb_i    :  IN STD_LOGIC;
         cp_i    :  IN STD_LOGIC;
          d_i    :  IN STD_LOGIC_VECTOR(87 DOWNTO 0);
         dv_i    :  IN STD_LOGIC;
         br_i    :  IN STD_LOGIC;
        txd_o    : OUT STD_LOGIC;
        trg_o    : OUT STD_LOGIC);
  END uat;
-- --------------------------------------------------------------------
   
