library IEEE;
use IEEE.STD_LOGIC_1164.ALL;
------------------------------------------------------------------------------------------------------------------------------
ENTITY TB_top_level IS	
END TB_top_level;
------------------------------------------------------------------------------------------------------------------------------
