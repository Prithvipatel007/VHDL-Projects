LIBRARY IEEE;
USE IEEE.STD_LOGIC_1164.ALL;
------------------------------------------------------------------------------------------------------------------------------
ENTITY brd_generator_e IS PORT(
    rb_i, cp_i, sel_i               :  IN STD_LOGIC;
    brd_o, clk_1k_o ,sec_o, secp_o  :  OUT STD_LOGIC
);
END brd_generator_e;
-------------------------------------------------------------------------------------------------------------------------------
