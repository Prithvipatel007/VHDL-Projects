library ieee;
use ieee.std_logic_1164.all;

entity tb_signal_generator_e is
end tb_signal_generator_e;