-- ----------------------------------------------------------------------------
-- ----------------------------------------------------------------------------
-- THIS FILE: sr08e_e.vhd - last edited: 2021-1202
-- ----------------------------------------------------------------------------
-- sr08e, 8-Bit-Shift-Register
-- ----------------------------------------------------------------------------
-- ----------------------------------------------------------------------------
  LIBRARY IEEE;
  USE IEEE.STD_LOGIC_1164.ALL;
--USE WORK.ifx_pack.ALL;
-- ----------------------------------------------------------------------------
  ENTITY sr08e IS
  PORT (rb_i,cp_i :  IN STD_LOGIC;
        en_i      :  IN STD_LOGIC;
        sdi_i     :  IN STD_LOGIC;
        q_o       : OUT STD_LOGIC_VECTOR (7 DOWNTO 0) );
  END sr08e;
-- ----------------------------------------------------------------------------
-- ----------------------------------------------------------------------------




