library ieee;
use ieee.std_logic_1164.all;

entity tb_morse_ascii_e is 
end tb_morse_ascii_e;

