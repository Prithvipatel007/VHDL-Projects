LIBRARY IEEE;
USE IEEE.STD_LOGIC_1164.ALL;

ENTITY tb_top_level_transmission_e IS
END tb_top_level_transmission_e;