library ieee;
use ieee.std_logic_1164.all;

entity tb_transmission_e is
end tb_transmission_e;