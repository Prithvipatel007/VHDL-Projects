LIBRARY IEEE;
USE IEEE.STD_LOGIC_1164.ALL;
-----------------------------------------------------------
ENTITY tb_shaper_e IS 
END tb_shaper_e;

