LIBRARY IEEE;
USE IEEE.STD_LOGIC_1164.ALL;
-----------------------------------------------------------------------------------------
ENTITY tb_tsc_ctrl_e IS END tb_tsc_ctrl_e;
--
