-- --------------------------------------------------------------------
-- --------------------------------------------------------------------
-- file: reg08_e.vhd, last modified: 2021-1202
-- --------------------------------------------------------------------
-- --------------------------------------------------------------------
-- some GHDL-cmds:   ghdl -s xxx.vhd  : Syntax check
--                   ghdl -a xxx.vhd  : Assembles file xxx.vhd
--                   ghdl -e xyz      : Elaborates xyz
-- prepare waveform: ghdl -r xxx_TB1 --wave=xxx_TB1_wave.ghw
-- --------------------------------------------------------------------
-- --------------------------------------------------------------------
  LIBRARY IEEE;
  USE IEEE.STD_LOGIC_1164.ALL;

  ENTITY reg08 IS    -- 8-bit-input-register 
   PORT (rb_i,cp_i  :  IN STD_LOGIC;
         en_i       :  IN STD_LOGIC;   -- enable to store data
         d_i        :  IN STD_LOGIC_VECTOR(7 DOWNTO 0);
         q_o        : OUT STD_LOGIC_VECTOR(7 DOWNTO 0) );
  END reg08;
--
-- ------------------------------------------------------------
-- ------------------------------------------------------------

