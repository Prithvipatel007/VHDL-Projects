-- --------------------------------------------------------------------
-- --------------------------------------------------------------------
-- THIS FILE: ifx_e.vhd - last edited: 2021-1202
-- --------------------------------------------------------------------
-- --------------------------------------------------------------------
-- ifx- The Serial Input Section
-- --------------------------------------------------------------------
-- --------------------------------------------------------------------
  LIBRARY IEEE;
  USE IEEE.STD_LOGIC_1164.ALL;
--USE WORK.ifx_pack.ALL;
-- --------------------------------------------------------------------
  ENTITY ifx IS
  PORT (rb_i   :  IN STD_LOGIC;                    -- Reset, active low
        cp_i   :  IN STD_LOGIC;                    -- Syscp, @ 12MHz
       sdi_i   :  IN STD_LOGIC;                    -- Serial Data 
       sdv_i   :  IN STD_LOGIC;                    -- Serial Data valid
       stx_i   :  IN STD_LOGIC;                    -- Transmitting now
         q_o   : OUT STD_LOGIC_VECTOR(87 DOWNTO 0);-- Data
        dv_o   : OUT STD_LOGIC);                   -- Data valid
  END ifx;
-- --------------------------------------------------------------------
-- --------------------------------------------------------------------


