LIBRARY IEEE;
USE IEEE.STD_LOGIC_1164.ALL;

ENTITY tb_morse_decoder_e IS 
END tb_morse_decoder_e;

