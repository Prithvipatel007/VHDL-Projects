library IEEE;
USE IEEE.STD_LOGIC_1164.ALL;

ENTITY TB_transmission_e IS 
END TB_transmission_e;

