LIBRARY IEEE;
USE IEEE.STD_LOGIC_1164.ALL;

ENTITY c10ec_e IS 
    PORT(
        rb_i,cp_i,en_i,cl_i     : IN STD_LOGIC;
        q3_o,co_o               : OUT STD_LOGIC);
END c10ec_e;

