library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;

entity tb_ascii_morse_e is
end tb_ascii_morse_e;