LIBRARY IEEE;
USE IEEE.STD_LOGIC_1164.ALL;

ENTITY tb_clock_divider_e IS
END tb_clock_divider_e;