library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;

entity tb_top_level_rx_e is
end tb_top_level_rx_e;