-- --------------------------------------------------------------------
-- --------------------------------------------------------------------
-- THIS FILE: c16ec_a1.vhd - last edited: 2021-1202
-- --------------------------------------------------------------------
-- --------------------------------------------------------------------
-- c10ec :  a 16-state-counter, has enable, has carry
-- --------------------------------------------------------------------
-- --------------------------------------------------------------------
-- some GHDL-cmds:   ghdl -s xxx.vhd  : Syntax check
--                   ghdl -a xxx.vhd  : Assembles file xxx.vhd
--                   ghdl -e xyz      : Elaborates xyz                
-- prepare waveform: ghdl -r xxx_TB1 --wave=xxx_TB1_wave.ghw
-- --------------------------------------------------------------------
-- --------------------------------------------------------------------
  LIBRARY IEEE;
  USE IEEE.STD_LOGIC_1164.ALL;
-- --------------------------------------------------------------------
  ENTITY c16ec IS   -- counter, mod10, has ena, has carry out
   PORT (rb_i,cp_i  :  IN STD_LOGIC;
         en_i       :  IN STD_LOGIC;                 -- enable counting
         co_o       : OUT STD_LOGIC);
  END c16ec;
-- --------------------------------------------------------------------

