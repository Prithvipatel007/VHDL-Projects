LIBRARY IEEE;
USE IEEE.STD_LOGIC_1164.ALL;
-----------------------------------------------------------------------------------------
ENTITY tb_gen_snd_e IS END tb_gen_snd_e;
--
