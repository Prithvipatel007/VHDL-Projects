-- --------------------------------------------------------------------
-- --------------------------------------------------------------------
-- THIS FILE: c05ec_a1.vhd - last edited: 2021-1202
-- --------------------------------------------------------------------
-- c05xc : a 5-state-counter, no enable, has carry
-- --------------------------------------------------------------------
-- --------------------------------------------------------------------
-- some GHDL-cmds:   ghdl -s xxx.vhd  : Syntax check
--                   ghdl -a xxx.vhd  : Assembles file xxx.vhd
--                   ghdl -e xyz      : Elaborates xyz
-- prepare waveform: ghdl -r xxx_TB1 --wave=xxx_TB1_wave.ghw
-- --------------------------------------------------------------------
-- --------------------------------------------------------------------
  LIBRARY IEEE;
  USE IEEE.STD_LOGIC_1164.ALL;
-- --------------------------------------------------------------------
-- counter, mod5, no ena, but carry out
--
  ENTITY c05xc IS   -- counter, mod5, no ena, but carry out
   PORT (rb_i,cp_i  :  IN STD_LOGIC;
         co_o       : OUT STD_LOGIC);
   END c05xc;
-- --------------------------------------------------------------------
-- --------------------------------------------------------------------

