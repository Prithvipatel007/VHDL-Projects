LIBRARY IEEE;
USE IEEE.STD_LOGIC_1164.ALL;
-----------------------------------------------------------------------------------------
ENTITY tb_ata_ctrl_e IS END tb_ata_ctrl_e;
--
