-- ----------------------------------------------------------------------------
-- ----------------------------------------------------------------------------
-- THIS FILE: sr08e_a1.vhd - last edited: 2021-1202
-- ----------------------------------------------------------------------------
-- ifx- The Serial Input Section, 8-Bit-Shift-Register
-- ----------------------------------------------------------------------------
-- --------------------------------------------------------------------
  LIBRARY IEEE;
  USE IEEE.STD_LOGIC_1164.ALL;
--USE WORK.ifx_pack.ALL;
-- --------------------------------------------------------------------
-- --------------------------------------------------------------------
-- shift sdi to q_o(7), q_o(7) to q_o(6),..., q_o(1) to q_o(0)
-- -------------------------------------------------------------------- 
  ARCHITECTURE a1 OF sr08e IS

  SIGNAL state_s : STD_LOGIC_VECTOR (7 DOWNTO 0);
-- -------------------------------------------------------------------- 
  BEGIN
  srx : PROCESS (rb_i,cp_i,state_s)
   BEGIN
   IF (rb_i='0') THEN state_s <= "00000000";
   ELSIF (cp_i='1' AND cp_i'EVENT)
    THEN
     IF  (en_i='1') THEN state_s(7)<=sdi_i;
                         state_s(6)<=state_s(7);
                         state_s(5)<=state_s(6);
                         state_s(4)<=state_s(5);
                         state_s(3)<=state_s(4);
                         state_s(2)<=state_s(3);
                         state_s(1)<=state_s(2);
                         state_s(0)<=state_s(1);
     END IF;
   END IF;
   END PROCESS srx;
-- -------------------------------------------------------------------- 
	q_o <= state_s;
-- -------------------------------------------------------------------- 
  END a1;
-- --------------------------------------------------------------------
